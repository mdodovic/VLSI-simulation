module testbench;

endmodule
