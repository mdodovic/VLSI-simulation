module testbench;


endmodule
