module m21_gate (
    I0,
    I1,
    S0,
    Y
);

    input I0, I1, S0;
    output Y;
    
endmodule