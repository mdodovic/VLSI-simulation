module helloWorldModule;

	initial begin
		$display("Hello world");
		$finish;
	end

endmodule
