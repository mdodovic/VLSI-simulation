module dut(clk, rst_n, t, q);

	input clk, rst_n, t;
	output q;

endmodule
