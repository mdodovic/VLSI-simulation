module testbench;
	
endmodule