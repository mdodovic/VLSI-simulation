module helloworld;

	initial begin
		$display("Hello world"); 
		$finish;		
	end

endmodule
